
-- Package for the use
package Register_pkg is
  
  -- Pulse for bit in register
  TYPE Pulse_State_Type IS (IDLE,PULSE,RESET);  -- Define the states
	
end Register_pkg;

package body Register_pkg is

end Register_pkg;
